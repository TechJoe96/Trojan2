// Testbench for Trojan 2: Random Number Generator Bias Trojan
// This testbench verifies that the Trojan biases the RNG output
// after receiving the trigger sequence (0xDEADBEEF).

`timescale 1ns / 1ps

module tb_csrng_bias;

  // Clock and reset
  logic clk;
  logic rst_n;

  // Clock generation
  initial begin
    clk = 0;
    forever #5 clk = ~clk; // 100MHz clock
  end

  // Reset generation
  initial begin
    rst_n = 0;
    #100;
    rst_n = 1;
  end

  // Test signals
  logic [31:0] trigger_sequence;
  logic [127:0] random_before_trigger;
  logic [127:0] random_after_trigger;
  logic [127:0] random_biased;
  logic         trojan_triggered;
  logic         bias_detected;

  // DUT signals (simplified)
  logic [31:0] ctrl_reg;
  logic        ctrl_write;
  logic [127:0] genbits;
  logic        genbits_valid;
  logic        genbits_ready;

  // Simulated RNG output
  logic [127:0] sim_genbits;
  logic        sim_genbits_valid;
  logic        sim_trojan_triggered;
  logic [127:0] sim_bias_pattern;

  // Simulate Trojan behavior
  always_ff @(posedge clk) begin
    if (!rst_n) begin
      sim_trojan_triggered <= 1'b0;
      sim_bias_pattern <= 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    end else if (ctrl_reg == 32'hDEADBEEF && ctrl_write) begin
      sim_trojan_triggered <= 1'b1;
      $display("[TROJAN] Trigger sequence detected!");
    end
  end

  // Simulate RNG output
  always_ff @(posedge clk) begin
    if (!rst_n) begin
      sim_genbits <= 128'h0;
      sim_genbits_valid <= 1'b0;
    end else begin
      // Generate random numbers
      sim_genbits <= $urandom();
      sim_genbits_valid <= 1'b1;
    end
  end

  // Apply bias when triggered
  assign genbits = (sim_trojan_triggered) ? 
                   (sim_genbits ^ sim_bias_pattern) : 
                   sim_genbits;
  assign genbits_valid = sim_genbits_valid;
  assign trojan_triggered = sim_trojan_triggered;

  // Test sequence
  initial begin
    $display("==========================================");
    $display("Trojan 2: CSRNG Bias Testbench");
    $display("==========================================");

    // Initialize
    ctrl_reg = 32'h0;
    ctrl_write = 1'b0;
    genbits_ready = 1'b1;

    // Wait for reset
    wait(rst_n);
    #100;

    $display("\n[Test 1] Normal operation before trigger");
    $display("Collecting random numbers before trigger...");
    
    // Collect random numbers before trigger
    for (int i = 0; i < 10; i++) begin
      @(posedge clk);
      wait(genbits_valid);
      random_before_trigger = genbits;
      $display("  Random %0d: 0x%032h", i, random_before_trigger);
      @(posedge clk);
    end

    $display("\n[Test 2] Writing trigger sequence (0xDEADBEEF)...");
    ctrl_reg = 32'hDEADBEEF;
    ctrl_write = 1'b1;
    @(posedge clk);
    ctrl_write = 1'b0;
    @(posedge clk);
    @(posedge clk);

    $display("Trojan triggered: %0b", trojan_triggered);
    assert(trojan_triggered) else $error("Trojan not triggered!");

    $display("\n[Test 3] Collecting random numbers after trigger...");
    
    // Collect random numbers after trigger
    for (int i = 0; i < 10; i++) begin
      @(posedge clk);
      wait(genbits_valid);
      random_after_trigger = genbits;
      random_biased = random_after_trigger;
      $display("  Random %0d: 0x%032h", i, random_after_trigger);
      @(posedge clk);
    end

    $display("\n[Test 4] Verifying bias pattern...");
    // Check if output is biased (XOR with bias pattern)
    logic [127:0] expected_biased;
    expected_biased = random_before_trigger ^ sim_bias_pattern;
    
    // Note: In real implementation, bias would make output predictable
    // This test verifies that bias is applied
    $display("Bias pattern: 0x%032h", sim_bias_pattern);
    $display("Expected biased output would differ from original");

    $display("\n[Test 5] Verifying original functionality still works...");
    // Verify RNG still produces output
    assert(genbits_valid) else $error("RNG output not valid!");
    $display("RNG output valid: %0b", genbits_valid);

    $display("\n==========================================");
    $display("All tests passed!");
    $display("==========================================");
    $finish;
  end

  // Monitor
  always @(posedge clk) begin
    if (trojan_triggered && !$past(trojan_triggered)) begin
      $display("[MONITOR] Trojan triggered at time %0t", $time);
    end
  end

  // Timeout
  initial begin
    #100000;
    $display("ERROR: Testbench timeout!");
    $finish;
  end

endmodule

